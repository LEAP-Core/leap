
import soft_connections::*;

import traffic_light_function::*;


module [CONNECTED_MODULE] mkSystem ();

   let tl <- mk_traffic_light();
  
endmodule
