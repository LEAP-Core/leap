../basic/channelio-common.bsv