`include "awb/provides/soft_connections.bsh"

`include "awb/provides/virtual_devices.bsh"


module [CONNECTED_MODULE] mkCommonServices#(VIRTUAL_DEVICES vdevs)
    // interface:
        ();

endmodule
