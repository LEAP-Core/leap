
`include "awb/provides/virtual_devices.bsh"

module mkStarterService#(VIRTUAL_DEVICES vdevs)
    // interface:
        ();
    
endmodule
