
import soft_connections::*;

`include "asim/provides/clock_test.bsh"


module [CONNECTED_MODULE] mkConnectedApplication ();

   let tl <- mkClockTest();
  
endmodule
