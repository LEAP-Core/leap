`include "awb/provides/central_cache_service.bsh"
`include "awb/provides/scratchpad_memory_service.bsh"
`include "awb/provides/shared_memory_service.bsh"
`include "awb/provides/librl_bsv_base.bsh"

`include "awb/provides/virtual_devices.bsh"
`include "awb/provides/soft_connections.bsh"


module [CONNECTED_MODULE] mkMemServices
    // interface:
        ();
    
    let centralCacheService     <- mkCentralCacheService();
    let scratchpadMemoryService <- mkScratchpadMemoryService(centralCacheService);
    let sharedMemoryService     <- mkSharedMemoryService();
    
endmodule
