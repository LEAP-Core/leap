//
// Copyright (C) 2009 Intel Corporation
//
// This program is free software; you can redistribute it and/or
// modify it under the terms of the GNU General Public License
// as published by the Free Software Foundation; either version 2
// of the License, or (at your option) any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program; if not, write to the Free Software
// Foundation, Inc., 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.
//

`include "asim/provides/soft_connections.bsh"

`include "asim/provides/streams.bsh"
`include "asim/provides/assertions_controller.bsh"
`include "asim/provides/params_controller.bsh"


interface CENTRAL_CONTROLLERS;
    interface ASSERTIONS_CONTROLLER assertsController;
    interface PARAMS_CONTROLLER paramsController;
endinterface

// ================ Standard Controller ===============

module [CONNECTED_MODULE] mkCentralControllers
    // interface:
    (CENTRAL_CONTROLLERS);

    // instantiate sub-controllers
    ASSERTIONS_CONTROLLER assertsCtrl <- mkAssertionsController();
    PARAMS_CONTROLLER     paramsCtrl  <- mkParamsController();

    interface assertsController = assertsCtrl;
    interface paramsController  = paramsCtrl;
endmodule
