`include "asim/provides/virtual_platform.bsh"

module mkApplication#(VIRTUAL_PLATFORM vp) ();

endmodule

