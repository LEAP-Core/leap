//
// Copyright (c) 2015, Intel Corporation
// All rights reserved.
//
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// Redistributions of source code must retain the above copyright notice, this
// list of conditions and the following disclaimer.
//
// Redistributions in binary form must reproduce the above copyright notice,
// this list of conditions and the following disclaimer in the documentation
// and/or other materials provided with the distribution.
//
// Neither the name of the Intel Corporation nor the names of its contributors
// may be used to endorse or promote products derived from this software
// without specific prior written permission.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
// ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT OWNER OR CONTRIBUTORS BE
// LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
// CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
// SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
// INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
// CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
// ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
// POSSIBILITY OF SUCH DAMAGE.
//

/**
 * @file rrr-debug-definitions.bsv
 * @author Kermin Fleming
 * @brief Defines typeclasses for RRR debuggers.
 */

`include "asim/provides/umf.bsh"

//  A typeclass for RRR debuggers. Each RRR entity has a different
//  type (by design), but a common debug interface. This typeclass 
//  allows us to write common debug infrastructure for each.

interface RRR_SERVER_DEBUG; 

    method Bool                                   notEmpty();
    method RRR_DEMARSHALLER_STATE                 demarshallerState();
    method UMF_METHOD_ID                          methodID();
    method UMF_SERVICE_ID                         serviceID();
    method UMF_PHY_CHANNEL_PVT                    sequenceNumber();
    method UMF_PHY_CHANNEL_PVT                    sequenceNumberLast();
    method Tuple3#(Bit#(64), Bit#(64), UMF_CHUNK) chunk();
    method Bool                                   misroutedPacket();
    method Bool                                   illegalMethod();
    method Bool                                   incorrectLength();
    method Bit#(64)                               totalPackets();
    method Bit#(64)                               totalChunks();
    method String                                 serviceName();

endinterface
