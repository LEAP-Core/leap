
module mkSharedMemoryService
    // interface:
        (Empty);
  messageM("Not Here?");    
endmodule
