//
// Copyright (c) 2014, Intel Corporation
// All rights reserved.
//
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// Redistributions of source code must retain the above copyright notice, this
// list of conditions and the following disclaimer.
//
// Redistributions in binary form must reproduce the above copyright notice,
// this list of conditions and the following disclaimer in the documentation
// and/or other materials provided with the distribution.
//
// Neither the name of the Intel Corporation nor the names of its contributors
// may be used to endorse or promote products derived from this software
// without specific prior written permission.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
// ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT OWNER OR CONTRIBUTORS BE
// LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
// CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
// SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
// INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
// CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
// ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
// POSSIBILITY OF SUCH DAMAGE.
//

import Clocks::*;
import ModuleContext::*;

`include "awb/provides/fpga_components.bsh"
`include "awb/provides/clocks_device.bsh"
`include "awb/provides/soft_services_lib.bsh"
`include "awb/provides/soft_services.bsh"
`include "awb/provides/soft_clocks_lib.bsh"

instance SOFT_SERVICE#(LOGICAL_CLOCK_INFO);

    module initializeServiceContext (LOGICAL_CLOCK_INFO);

        let clock <- exposeCurrentClock();
        let reset <- exposeCurrentReset();

        return LOGICAL_CLOCK_INFO {clk: clock, rst: reset};

    endmodule
    
    module finalizeServiceContext#(LOGICAL_CLOCK_INFO info) (Empty);
        // Currently nothing to do here.
    endmodule

endinstance

instance SYNTHESIZABLE_SOFT_SERVICE#(LOGICAL_CLOCK_INFO, Empty);

    module exposeServiceContext#(LOGICAL_CLOCK_INFO info) (Empty);
        // Currently nothing to do here.
    endmodule

endinstance


module [t_CONTEXT] mkSoftClock#(Integer outputFreq) (UserClock)
    provisos
        (Context#(t_CONTEXT, LOGICAL_CLOCK_INFO),
         IsModule#(t_CONTEXT, t_DUMMY));

   // Get a reference to the known clock
   LOGICAL_CLOCK_INFO modelClock <- getContext();
   let returnClock <- mkUserClockFromFrequency(`MODEL_CLOCK_FREQ,
                                               outputFreq,
                                               clocked_by modelClock.clk, 
                                               reset_by modelClock.rst);
   return returnClock;
endmodule
