
typedef enum {
  Filling,
  Draining
} State deriving (Bits,Eq);

