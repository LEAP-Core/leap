import hasim_common::*;
import afu_alg::*;

module [HASIM_MODULE] mkSystem ();
   
  let alg <- mkAFU_Alg();
  
endmodule
