//
// Copyright (c) 2014, Intel Corporation
// All rights reserved.
//
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// Redistributions of source code must retain the above copyright notice, this
// list of conditions and the following disclaimer.
//
// Redistributions in binary form must reproduce the above copyright notice,
// this list of conditions and the following disclaimer in the documentation
// and/or other materials provided with the distribution.
//
// Neither the name of the Intel Corporation nor the names of its contributors
// may be used to endorse or promote products derived from this software
// without specific prior written permission.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
// ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT OWNER OR CONTRIBUTORS BE
// LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
// CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
// SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
// INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
// CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
// ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
// POSSIBILITY OF SUCH DAMAGE.
//

`include "awb/provides/low_level_platform_interface.bsh"

`include "awb/rrr/client_stub_STARTER_DEVICE.bsh"
`include "awb/rrr/server_stub_STARTER_DEVICE.bsh"

// Starter
interface STARTER;

    // server methods
    method Action acceptRequest_Start();

    // client methods
    method Action makeRequest_End(Bit#(8) exit_code);
    
    //
    // FPGA Heartbeat --
    //   Message the number of FPGA cycles passed.
    //   Useful for detecting deadlocks.
    //
    method Action makeRequest_Heartbeat(Bit#(64) fpga_cycles);

endinterface

// mkStarter
module [CONNECTED_MODULE] mkStarter#(LowLevelPlatformInterface llpi)
    // interface:
        (STARTER);

    // ----------- stubs -----------
    ClientStub_STARTER_DEVICE client_stub <- mkClientStub_STARTER_DEVICE;
    ServerStub_STARTER_DEVICE server_stub <- mkServerStub_STARTER_DEVICE;
    
    // ----------- server methods ------------

    // Run
    method Action acceptRequest_Start ();
        let r <- server_stub.acceptRequest_Start();
    endmethod

    // ------------ client methods ------------

    // signal end of simulation
    method Action makeRequest_End(Bit#(8) exit_code);
        client_stub.makeRequest_End(exit_code);
    endmethod

    // Heartbeat
    method Action makeRequest_Heartbeat(Bit#(64) fpga_cycles);
        client_stub.makeRequest_Heartbeat(fpga_cycles);
    endmethod

endmodule
