import hasim_common::*;
import dme_alg::*;

module [HASIM_MODULE] mkSystem ();
   
  let alg <- mkDME_Alg();
  
endmodule
