// Need to include some stuff here. 
//`include "soft_services.bsv"