
`include "awb/provides/virtual_devices.bsh"
`include "awb/provides/shared_memory.bsh"

`include "awb/provides/soft_connections.bsh"


module [CONNECTED_MODULE] mkSharedMemoryService#(VIRTUAL_DEVICES vdevs)
    // interface:
        (Empty);
  messageM("Not Here?");    
endmodule
