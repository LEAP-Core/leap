`include "hasim_common.bsh"

//=============== Null Controller ===============
module [HASIM_MODULE] mkController();
endmodule

