// Need to include some stuff here. 