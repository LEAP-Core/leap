`include "asim/provides/fpga_components.bsh"
`include "asim/provides/clocks_device.bsh"
// Need the lib seperation to prevent death by AWB

typedef UserClock LOGICAL_CLOCK_INFO;




