
`include "awb/provides/virtual_devices.bsh"


module mkFrontPanelService#(VIRTUAL_DEVICES vdevs)
    // interface:
        ();

endmodule
