`include "asim/provides/soft_connections.bsh"

`include "asim/provides/traffic_light_function.bsh"


module [CONNECTED_MODULE] mkSystem ();

  let tl <- mkTrafficLightFunction();

endmodule
